`timescale 1ns / 1ps

module spare_allocation_analyzer (
	input 
);


endmodule