`timescale 1ns / 1ps

module RedundantAnalyzer (
	input [4:0] unused_spare,
	input uncover_must_pivot,
	input signal_valid,
	input [PCAM-1:0][4:0] uncover_nonpivot_addr,
	input [4:0] cover_pivot_addr [0:4],
	input [7:0] nonpivot_cover_result,
	input uncover_must_addr,
	output final_result,
	output [15:0] final_cover_addr
);

parameter PCAM = 8;
parameter NPCAM = 30;



<<<<<<<< HEAD:Verilog/RedundantAnalyzer.v


========
>>>>>>>> f0f68ffc7309aba7898667a811948d61414a1cc7:Verilog/redundant_analyzer.v
endmodule
